module SB_HFOSC;
endmodule

module SB_PLL40_CORE;
endmodule


